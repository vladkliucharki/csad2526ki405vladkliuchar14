/*
 * Module: i2c_master_rx (I2C Master Receiver / Decoder)
 * Language: Verilog
 * Task: 14
 *
 * Purpose: 
 * Implements I2C Master logic for receiving one byte of data (Read).
 * Generates clock pulses (SCL) and controls the data flow (SDA).
 */
module i2c_master_rx (
    // --- System Ports ---
    input wire           clk,        // System clock signal
    input wire           rst_n,      // Asynchronous active-low reset

    // --- User Control Ports ---
    input wire           start_rx,   // Pulse to start transaction
    input wire [6:0]     slave_addr, // 7-bit Slave device address

    // --- Status and Data Ports ---
    output wire          busy,       // '1' - transaction in progress
    output wire          ack_error,  // '1' - if NACK is received (error)
    output wire [7:0]    data_out,   // 8-bit received data byte
    output wire          data_ready  // '1' - pulse, data_out is valid

    // --- I2C Bus Ports ---
    inout wire           sda,        // Bidirectional I2C data line
    output wire          scl         // I2C clock line (generated by master)
);

    // =========================================================================
    // --- Clock Divider Parameters ---
    // =========================================================================
    parameter CLK_FREQ = 50_000_000;
    parameter I2C_FREQ = 100_000;
    localparam HALF_PERIOD_COUNT = (CLK_FREQ / (I2C_FREQ * 2)) - 1;

    // =========================================================================
    // --- Internal Registers and Signals ---
    // =========================================================================
    
    // --- Clock Divider ---
    reg [$clog2(HALF_PERIOD_COUNT):0] clk_div_cnt;
    reg tick;

    // --- FSM Registers ---
    reg [4:0] state;
    reg busy_reg;
    reg ack_error_reg;
    reg data_ready_reg;
    
    // --- Bus Control Registers ---
    reg scl_reg;
    reg sda_o_reg;
    reg sda_en_reg;

    // --- Data Registers ---
    reg [7:0] shift_reg;   // Shift register (for address + R/W, and data reception)
    reg [7:0] data_out_reg;
    reg [2:0] bit_cnt;

    // --- FSM States ---
    localparam S_IDLE             = 5'd0;  // Idle
    localparam S_START_1          = 5'd1;  // Generate START
    localparam S_START_2          = 5'd2;
    localparam S_TX_ADDR_BIT      = 5'd3;  // Transmit address bit
    localparam S_TX_ADDR_CLK_HI   = 5'd4;
    localparam S_TX_ADDR_CLK_LO   = 5'd5;
    localparam S_GET_ADDR_ACK_1   = 5'd6;  // Receive ACK (after address)
    localparam S_GET_ADDR_ACK_CLK = 5'd7;
    localparam S_GET_ADDR_ACK_RD  = 5'd8;
    localparam S_GET_ADDR_ACK_LO  = 5'd9;
    localparam S_RX_CLK_HI        = 5'd10; // Receive data bit
    localparam S_RX_BIT_READ      = 5'd11;
    localparam S_RX_CLK_LO        = 5'd12;
    localparam S_SEND_NACK_1      = 5'd13; // Send NACK (end of read)
    localparam S_SEND_NACK_CLK_HI = 5'd14;
    localparam S_SEND_NACK_CLK_LO = 5'd15;
    localparam S_STOP_1           = 5'd16; // Generate STOP
    localparam S_STOP_CLK_HI      = 5'd17;
    localparam S_STOP_2           = 5'd18;

    // =========================================================================
    // --- Output Assignments ---
    // =========================================================================
    assign scl = scl_reg;
    assign sda = (sda_en_reg) ? sda_o_reg : 1'bz;
    assign busy = busy_reg;
    assign ack_error = ack_error_reg;
    assign data_out = data_out_reg;
    assign data_ready = data_ready_reg;

    // =========================================================================
    // --- Clock Divider Logic ---
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            clk_div_cnt <= 0;
            tick <= 1'b0;
        end else begin
            if (clk_div_cnt == HALF_PERIOD_COUNT) begin
                clk_div_cnt <= 0;
                tick <= 1'b1;
            end else begin
                clk_div_cnt <= clk_div_cnt + 1;
                tick <= 1'b0;
            end
        end
    end

    // =========================================================================
    // --- FSM (Finite State Machine) Logic ---
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // Reset to initial state
            state <= S_IDLE;
            scl_reg <= 1'b1; sda_o_reg <= 1'b1; sda_en_reg <= 1'b1;
            busy_reg <= 1'b0; ack_error_reg <= 1'b0; data_ready_reg <= 1'b0;
            data_out_reg <= 0; bit_cnt <= 0; shift_reg <= 0;
            
        end else if (tick) begin 
            
            // data_ready is a pulse, reset it by default
            data_ready_reg <= 1'b0;
            
            case (state)
                
                // --- Idle State ---
                S_IDLE: begin
                    busy_reg <= 1'b0;
                    ack_error_reg <= 1'b0;
                    scl_reg <= 1'b1; sda_o_reg <= 1'b1; sda_en_reg <= 1'b1; 
                    
                    if (start_rx) begin
                        busy_reg <= 1'b1;
                        state <= S_START_1;
                    end
                end

                // --- START Condition ---
                S_START_1: begin
                    sda_o_reg <= 1'b0;
                    state <= S_START_2;
                end
                
                S_START_2: begin
                    scl_reg <= 1'b0;
                    // Load address and R/W=1 bit (Read)
                    shift_reg <= {slave_addr, 1'b1}; 
                    bit_cnt <= 3'd7; 
                    state <= S_TX_ADDR_BIT;
                end

                // --- Transmit Bit (Address) ---
                S_TX_ADDR_BIT: begin
                    sda_o_reg <= shift_reg[7];
                    state <= S_TX_ADDR_CLK_HI;
                end
                
                S_TX_ADDR_CLK_HI: begin
                    scl_reg <= 1'b1;
                    state <= S_TX_ADDR_CLK_LO;
                end
                
                S_TX_ADDR_CLK_LO: begin
                    scl_reg <= 1'b0;
                    if (bit_cnt == 0) begin
                        state <= S_GET_ADDR_ACK_1;
                    end else begin
                        shift_reg <= shift_reg << 1;
                        bit_cnt <= bit_cnt - 1;
                        state <= S_TX_ADDR_BIT;
                    end
                end

                // --- Receive ACK/NACK (after Address) ---
                S_GET_ADDR_ACK_1: begin
                    sda_en_reg <= 1'b0; // "Release" SDA
                    state <= S_GET_ADDR_ACK_CLK;
                end
                
                S_GET_ADDR_ACK_CLK: begin
                    scl_reg <= 1'b1;
                    state <= S_GET_ADDR_ACK_RD;
                end
                
                S_GET_ADDR_ACK_RD: begin
                    if (sda == 1'b1) begin // '1' == NACK
                        ack_error_reg <= 1'b1;
                    end
                    state <= S_GET_ADDR_ACK_LO;
                end

                S_GET_ADDR_ACK_LO: begin
                    scl_reg <= 1'b0;
                    if (ack_error_reg) begin
                        sda_en_reg <= 1'b1; // Regain control
                        state <= S_STOP_1;  // Error, stop
                    end else begin
                        // Received ACK, preparing to receive data
                        bit_cnt <= 3'd7; 
                        shift_reg <= 0;  // Clear shift register
                        state <= S_RX_CLK_HI;
                        // sda_en_reg remains '0' (Hi-Z) because we are listening
                    end
                end

                // --- Receive Data Byte ---
                S_RX_CLK_HI: begin
                    scl_reg <= 1'b1; // SCL=1
                    state <= S_RX_BIT_READ;
                end

                S_RX_BIT_READ: begin
                    // Read bit from SDA (while SCL=1)
                    shift_reg <= {shift_reg[6:0], sda}; // Shift and write
                    state <= S_RX_CLK_LO;
                end
                
                S_RX_CLK_LO: begin
                    scl_reg <= 1'b0; // SCL=0
                    if (bit_cnt == 0) begin
                        // Received all 8 bits
                        data_out_reg <= shift_reg; // Save the result
                        data_ready_reg <= 1'b1;    // Signal data ready
                        state <= S_SEND_NACK_1;    // Send NACK (end of reception)
                    end else begin
                        bit_cnt <= bit_cnt - 1;
                        state <= S_RX_CLK_HI; // Next bit
                    end
                end

                // --- Send NACK (end of read) ---
                S_SEND_NACK_1: begin
                    // We (Master) send NACK to tell the Slave "stop"
                    sda_en_reg <= 1'b1;    // Take control of SDA
                    sda_o_reg <= 1'b1;     // Set '1' (NACK)
                    state <= S_SEND_NACK_CLK_HI;
                end
                
                S_SEND_NACK_CLK_HI: begin
                    scl_reg <= 1'b1;
                    state <= S_SEND_NACK_CLK_LO;
                end
                
                S_SEND_NACK_CLK_LO: begin
                    scl_reg <= 1'b0;
                    state <= S_STOP_1; // Go to STOP
                end

                // --- STOP Condition ---
                S_STOP_1: begin
                    sda_en_reg <= 1'b1;
                    sda_o_reg <= 1'b0;
                    state <= S_STOP_CLK_HI;
                end

                S_STOP_CLK_HI: begin
                    scl_reg <= 1'b1;
                    state <= S_STOP_2;
                end
                
                S_STOP_2: begin
                    sda_o_reg <= 1'b1;
                    state <= S_IDLE;
                end
                
                default: begin
                    state <= S_IDLE;
                end
                
            endcase
        end
    end

endmodule