/*
 * Module: i2c_master_tx (I2C Master Transmitter / Encoder)
 * Language: Verilog
 * Task: 14
 *
 * Purpose: 
 * Implements I2C Master logic for transmitting one byte of data (Write).
 * Generates clock pulses (SCL) and controls the data flow (SDA).
 */
module i2c_master_tx (
    // --- System Ports ---
    input wire           clk,        // System clock signal (e.g., 50 MHz)
    input wire           rst_n,      // Asynchronous active-low reset

    // --- User Control Ports ---
    input wire           start_tx,   // Pulse to start transaction
    input wire [6:0]     slave_addr, // 7-bit Slave device address
    input wire [7:0]     data_in,    // 8-bit data byte for transmission

    // --- Status Ports ---
    output wire          busy,       // '1' - transaction in progress, '0' - ready
    output wire          ack_error,  // '1' - if NACK is received (error)

    // --- I2C Bus Ports ---
    inout wire           sda,        // Bidirectional I2C data line
    output wire          scl         // I2C clock line (generated by master)
);

    // =========================================================================
    // --- Clock Divider Parameters ---
    // =========================================================================
    // Set your system clock frequency
    parameter CLK_FREQ = 50_000_000;  // Example: 50 MHz
    // Desired SCL frequency (100 kHz for Standard Mode)
    parameter I2C_FREQ = 100_000;
    
    // Calculation of the divider to get *half* the SCL period.
    // The FSM (Finite State Machine) will operate on "ticks" at 2x I2C_FREQ.
    localparam HALF_PERIOD_COUNT = (CLK_FREQ / (I2C_FREQ * 2)) - 1;

    // =========================================================================
    // --- Internal Registers and Signals ---
    // =========================================================================
    
    // --- Clock Divider ---
    reg [$clog2(HALF_PERIOD_COUNT):0] clk_div_cnt; // Divider counter
    reg tick;                                      // Output "tick" for FSM

    // --- FSM (Finite State Machine) Registers ---
    reg [4:0] state;       // FSM current state register
    reg busy_reg;          // Internal 'busy' register
    reg ack_error_reg;     // Internal 'ack_error' register
    
    // --- Bus Control Registers ---
    reg scl_reg;           // Register for controlling scl output
    reg sda_o_reg;         // Register for the *value* of sda output
    reg sda_en_reg;        // Register for *enabling* sda output ('1' = output, '0' = input/Hi-Z)

    // --- Data Registers ---
    reg [7:0] shift_reg;   // Shift register (for address + R/W bit, and data)
    reg [2:0] bit_cnt;     // Bit counter (0-7)
    reg       sending_addr;  // '1' - sending address, '0' - sending data

    // --- FSM States ---
    localparam S_IDLE             = 5'd0;  // Idle
    localparam S_START_1          = 5'd1;  // Generate START: SDA=0 (SCL=1)
    localparam S_START_2          = 5'd2;  // Generate START: SCL=0
    localparam S_TX_BIT           = 5'd3;  // Set bit on SDA (SCL=0)
    localparam S_TX_CLK_HI        = 5'd4;  // SCL=1 (Slave reads bit)
    localparam S_TX_CLK_LO        = 5'd5;  // SCL=0 (End of bit transmission)
    localparam S_GET_ACK_1        = 5'd6;  // Release SDA (for ACK)
    localparam S_GET_ACK_CLK_HI   = 5'd7;  // SCL=1 (for ACK)
    localparam S_GET_ACK_READ     = 5'd8;  // Read ACK/NACK from SDA
    localparam S_GET_ACK_CLK_LO   = 5'd9;  // SCL=0 (for ACK)
    localparam S_STOP_1           = 5'd10; // Generate STOP: SDA=0 (SCL=0)
    localparam S_STOP_CLK_HI      = 5'd11; // Generate STOP: SCL=1
    localparam S_STOP_2           = 5'd12; // Generate STOP: SDA=1 (SCL=1)

    // =========================================================================
    // --- Output Assignments ---
    // =========================================================================
    
    // SCL Control: simply output the value from the register
    assign scl = scl_reg;
    
    // SDA Control: tri-state buffer.
    // sda_en_reg = 1 -> Master controls the line (outputs sda_o_reg).
    // sda_en_reg = 0 -> Master "releases" the line (Hi-Z), so Slave can send ACK.
    assign sda = (sda_en_reg) ? sda_o_reg : 1'bz;

    assign busy = busy_reg;
    assign ack_error = ack_error_reg;

    // =========================================================================
    // --- Clock Divider Logic ---
    // =========================================================================
    // Generates a 'tick' every HALF_PERIOD_COUNT 'clk' cycles.
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            clk_div_cnt <= 0;
            tick <= 1'b0;
        end else begin
            if (clk_div_cnt == HALF_PERIOD_COUNT) begin
                clk_div_cnt <= 0;
                tick <= 1'b1;
            end else begin
                clk_div_cnt <= clk_div_cnt + 1;
                tick <= 1'b0;
            end
        end
    end

    // =========================================================================
    // --- FSM (Finite State Machine) Logic ---
    // =========================================================================
    // All Master logic is implemented here.
    // Changes states only on 'tick'.
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // Reset to initial state
            state <= S_IDLE;
            scl_reg <= 1'b1;       // SCL "released" (high)
            sda_o_reg <= 1'b1;     // SDA "released" (high)
            sda_en_reg <= 1'b1;    // Driving the line
            busy_reg <= 1'b0;
            ack_error_reg <= 1'b0;
            bit_cnt <= 0;
            shift_reg <= 0;
            sending_addr <= 1'b0;
            
        end else if (tick) begin // Operate only on the "tick" from the divider
            
            case (state)
                
                // --- Idle State ---
                S_IDLE: begin
                    busy_reg <= 1'b0;
                    ack_error_reg <= 1'b0;
                    scl_reg <= 1'b1;
                    sda_o_reg <= 1'b1;
                    sda_en_reg <= 1'b1; 
                    
                    if (start_tx) begin
                        busy_reg <= 1'b1;
                        sending_addr <= 1'b1; // Start by sending the address
                        state <= S_START_1;
                    end
                end

                // --- START Condition ---
                S_START_1: begin
                    sda_o_reg <= 1'b0; // SCL=1, pull SDA=0
                    state <= S_START_2;
                end
                
                S_START_2: begin
                    scl_reg <= 1'b0; // Pull SCL=0. START condition generated.
                    // Load address and R/W=0 bit (Write)
                    shift_reg <= {slave_addr, 1'b0}; 
                    bit_cnt <= 3'd7; // We will transmit 8 bits
                    state <= S_TX_BIT;
                end

                // --- Bit Transmission ---
                S_TX_BIT: begin
                    sda_o_reg <= shift_reg[7]; // Set the MSB on SDA
                    state <= S_TX_CLK_HI;
                end
                
                S_TX_CLK_HI: begin
                    scl_reg <= 1'b1; // Raise SCL=1. Slave reads bit.
                    state <= S_TX_CLK_LO;
                end
                
                S_TX_CLK_LO: begin
                    scl_reg <= 1'b0; // Pull SCL=0.
                    if (bit_cnt == 0) begin
                        state <= S_GET_ACK_1; // 8 bits transmitted, wait for ACK
                    end else begin
                        shift_reg <= shift_reg << 1; // Shift the register
                        bit_cnt <= bit_cnt - 1;
                        state <= S_TX_BIT; // Next bit
                    end
                end

                // --- Receiving ACK/NACK ---
                S_GET_ACK_1: begin
                    sda_en_reg <= 1'b0; // "Release" SDA
                    state <= S_GET_ACK_CLK_HI;
                end
                
                S_GET_ACK_CLK_HI: begin
                    scl_reg <= 1'b1; // Clock SCL=1 for ACK
                    state <= S_GET_ACK_READ;
                end
                
                S_GET_ACK_READ: begin
                    if (sda == 1'b1) begin // '1' == NACK (error)
                        ack_error_reg <= 1'b1;
                    end
                    state <= S_GET_ACK_CLK_LO;
                end

                S_GET_ACK_CLK_LO: begin
                    scl_reg <= 1'b0; // Pull SCL=0
                    sda_en_reg <= 1'b1; // Regain control of SDA
                    
                    if (ack_error_reg) begin
                        state <= S_STOP_1; // Received NACK, stop
                    end else if (sending_addr) begin
                        // Received ACK after address, now send data
                        sending_addr <= 1'b0;
                        shift_reg <= data_in; // Load data
                        bit_cnt <= 3'd7;
                        state <= S_TX_BIT;
                    end else begin
                        // Received ACK after data, finish
                        state <= S_STOP_1;
                    end
                end

                // --- STOP Condition ---
                S_STOP_1: begin
                    sda_o_reg <= 1'b0; // SCL=0, SDA=0
                    state <= S_STOP_CLK_HI;
                end

                S_STOP_CLK_HI: begin
                    scl_reg <= 1'b1; // SCL=1
                    state <= S_STOP_2;
                end
                
                S_STOP_2: begin
                    sda_o_reg <= 1'b1; // SCL=1, SDA=1 -> STOP
                    state <= S_IDLE; // Return to idle
                end
                
                default: begin
                    state <= S_IDLE;
                end
                
            endcase
        end
    end

endmodule